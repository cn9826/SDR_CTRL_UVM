`define  APP_AW    26  // Application Address Width
`define  APP_DW    32  // Application Data Width 
`define  APP_BW    4  // Application Byte Width
`define  APP_RW    9  // Application Request Width

`define  SDR_DW    8 // SDR Data Width 
`define  SDR_BW    1   // SDR Byte Width

`define SDR_RFSH_TIMER_W 	12
`define SDR_RFSH_ROW_CNT_W	 3
